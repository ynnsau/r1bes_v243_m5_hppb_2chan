// (C) 2001-2024 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


// pcie_ed_pio0.v

// Generated using ACDS version 22.1 174

`timescale 1 ps / 1 ps
module pcie_ed_pio0 (
		input  wire          Clk_i,                    //              clk.clk
		input  wire          Rstn_i,                   //            reset.reset_n
		output wire          pio_clk,                  //   pio_master_clk.clk
		output wire          pio_rst_n,                // pio_master_reset.reset_n
		output wire [63:0]   pio_address_o,            //       pio_master.address
		output wire          pio_read_o,               //                 .read
		input  wire [1023:0] pio_readdata_i,           //                 .readdata
		input  wire          pio_readdatavalid_i,      //                 .readdatavalid
		output wire          pio_write_o,              //                 .write
		output wire [1023:0] pio_writedata_o,          //                 .writedata
		input  wire          pio_waitrequest_i,        //                 .waitrequest
		output wire [127:0]  pio_byteenable_o,         //                 .byteenable
		input  wire [1:0]    pio_response_i,           //                 .response
		output wire [3:0]    pio_burstcount_o,         //                 .burstcount
		input  wire [255:0]  pio_rx_st0_payload_i,     //       rx_st0_pio.data
		input  wire          pio_rx_st0_sop_i,         //                 .startofpacket
		input  wire          pio_rx_st0_eop_i,         //                 .endofpacket
		input  wire          pio_rx_st0_dvalid_i,      //                 .valid
		input  wire [2:0]    pio_rx_st0_empty_i,       //                 .empty
		output wire          pio_rx_st_ready_o,        //                 .ready
		input  wire [255:0]  pio_rx_st1_payload_i,     //       rx_st1_pio.data
		input  wire          pio_rx_st1_sop_i,         //                 .startofpacket
		input  wire          pio_rx_st1_eop_i,         //                 .endofpacket
		input  wire          pio_rx_st1_dvalid_i,      //                 .valid
		input  wire [2:0]    pio_rx_st1_empty_i,       //                 .empty
		input  wire [255:0]  pio_rx_st2_payload_i,     //       rx_st2_pio.data
		input  wire          pio_rx_st2_sop_i,         //                 .startofpacket
		input  wire          pio_rx_st2_eop_i,         //                 .endofpacket
		input  wire          pio_rx_st2_dvalid_i,      //                 .valid
		input  wire [2:0]    pio_rx_st2_empty_i,       //                 .empty
		input  wire [255:0]  pio_rx_st3_payload_i,     //       rx_st3_pio.data
		input  wire          pio_rx_st3_sop_i,         //                 .startofpacket
		input  wire          pio_rx_st3_eop_i,         //                 .endofpacket
		input  wire          pio_rx_st3_dvalid_i,      //                 .valid
		input  wire [2:0]    pio_rx_st3_empty_i,       //                 .empty
		output wire [2:0]    rx_st_hcrdt_init_o,       //  rx_st0_pio_misc.rx_st_Hcrdt_init
		output wire [2:0]    rx_st_hcrdt_update_o,     //                 .rx_st_Hcrdt_update
		output wire [5:0]    rx_st_hcrdt_update_cnt_o, //                 .rx_st_Hcrdt_update_cnt
		input  wire [2:0]    rx_st_hcrdt_init_ack_i,   //                 .rx_st_Hcrdt_init_ack
		output wire [2:0]    rx_st_dcrdt_init_o,       //                 .rx_st_Dcrdt_init
		output wire [2:0]    rx_st_dcrdt_update_o,     //                 .rx_st_Dcrdt_update
		output wire [11:0]   rx_st_dcrdt_update_cnt_o, //                 .rx_st_Dcrdt_update_cnt
		input  wire [2:0]    rx_st_dcrdt_init_ack_i,   //                 .rx_st_Dcrdt_init_ack
		input  wire [127:0]  pio_rx_st0_header_i,      //                 .rx_st0_hdr
		input  wire [31:0]   pio_rx_st0_tlp_prfx_i,    //                 .rx_st0_prefix
		input  wire          pio_rx_st0_hvalid_i,      //                 .rx_st0_hvalid
		input  wire          pio_rx_st0_pvalid_i,      //                 .rx_st0_pvalid
		input  wire [2:0]    pio_rx_st0_bar_i,         //                 .rx_st0_bar
		input  wire [127:0]  pio_rx_st1_header_i,      //                 .rx_st1_hdr
		input  wire [31:0]   pio_rx_st1_tlp_prfx_i,    //                 .rx_st1_prefix
		input  wire          pio_rx_st1_hvalid_i,      //                 .rx_st1_hvalid
		input  wire          pio_rx_st1_pvalid_i,      //                 .rx_st1_pvalid
		input  wire [2:0]    pio_rx_st1_bar_i,         //                 .rx_st1_bar
		input  wire [127:0]  pio_rx_st2_header_i,      //                 .rx_st2_hdr
		input  wire [31:0]   pio_rx_st2_tlp_prfx_i,    //                 .rx_st2_prefix
		input  wire          pio_rx_st2_hvalid_i,      //                 .rx_st2_hvalid
		input  wire          pio_rx_st2_pvalid_i,      //                 .rx_st2_pvalid
		input  wire [2:0]    pio_rx_st2_bar_i,         //                 .rx_st2_bar
		input  wire [127:0]  pio_rx_st3_header_i,      //                 .rx_st3_hdr
		input  wire [31:0]   pio_rx_st3_tlp_prfx_i,    //                 .rx_st3_prefix
		input  wire          pio_rx_st3_hvalid_i,      //                 .rx_st3_hvalid
		input  wire          pio_rx_st3_pvalid_i,      //                 .rx_st3_pvalid
		input  wire [2:0]    pio_rx_st3_bar_i,         //                 .rx_st3_bar
		output wire [255:0]  pio_tx_st0_payload_o,     //       tx_st0_pio.data
		output wire          pio_tx_st0_sop_o,         //                 .startofpacket
		output wire          pio_tx_st0_eop_o,         //                 .endofpacket
		output wire          pio_tx_st0_dvalid_o,      //                 .valid
		input  wire          pio_tx_st_ready_i,        //                 .ready
		output wire [255:0]  pio_tx_st1_payload_o,     //       tx_st1_pio.data
		output wire          pio_tx_st1_sop_o,         //                 .startofpacket
		output wire          pio_tx_st1_eop_o,         //                 .endofpacket
		output wire          pio_tx_st1_dvalid_o,      //                 .valid
		output wire [255:0]  pio_tx_st2_payload_o,     //       tx_st2_pio.data
		output wire          pio_tx_st2_sop_o,         //                 .startofpacket
		output wire          pio_tx_st2_eop_o,         //                 .endofpacket
		output wire          pio_tx_st2_dvalid_o,      //                 .valid
		output wire [255:0]  pio_tx_st3_payload_o,     //       tx_st3_pio.data
		output wire          pio_tx_st3_sop_o,         //                 .startofpacket
		output wire          pio_tx_st3_eop_o,         //                 .endofpacket
		output wire          pio_tx_st3_dvalid_o,      //                 .valid
		output wire [127:0]  pio_tx_st0_header_o,      //  tx_st0_pio_misc.tx_st0_hdr
		output wire [127:0]  pio_tx_st1_header_o,      //                 .tx_st1_hdr
		output wire [127:0]  pio_tx_st2_header_o,      //                 .tx_st2_hdr
		output wire [127:0]  pio_tx_st3_header_o,      //                 .tx_st3_hdr
		input  wire [2:0]    tx_st_hcrdt_init_i,       //                 .tx_st_Hcrdt_init
		input  wire [2:0]    tx_st_hcrdt_update_i,     //                 .tx_st_Hcrdt_update
		input  wire [5:0]    tx_st_hcrdt_update_cnt_i, //                 .tx_st_Hcrdt_update_cnt
		output wire [2:0]    tx_st_hcrdt_init_ack_o,   //                 .tx_st_Hcrdtt_init_ack
		input  wire [2:0]    tx_st_dcrdt_init_i,       //                 .tx_st_Dcrdt_init
		input  wire [2:0]    tx_st_dcrdt_update_i,     //                 .tx_st_Dcrdt_update
		input  wire [11:0]   tx_st_dcrdt_update_cnt_i, //                 .tx_st_Dcrdt_update_cnt
		output wire [2:0]    tx_st_dcrdt_init_ack_o,   //                 .tx_st_Dcrdt_init_ack
		output wire [31:0]   pio_tx_st0_prefix_o,      //                 .tx_st0_prefix
		output wire          pio_tx_st0_hvalid_o,      //                 .tx_st0_hvalid
		output wire          pio_tx_st0_pvalid_o,      //                 .tx_st0_pvalid
		output wire [31:0]   pio_tx_st1_prefix_o,      //                 .tx_st1_prefix
		output wire          pio_tx_st1_hvalid_o,      //                 .tx_st1_hvalid
		output wire          pio_tx_st1_pvalid_o,      //                 .tx_st1_pvalid
		output wire [31:0]   pio_tx_st2_prefix_o,      //                 .tx_st2_prefix
		output wire          pio_tx_st2_hvalid_o,      //                 .tx_st2_hvalid
		output wire          pio_tx_st2_pvalid_o,      //                 .tx_st2_pvalid
		output wire [31:0]   pio_tx_st3_prefix_o,      //                 .tx_st3_prefix
		output wire          pio_tx_st3_hvalid_o,      //                 .tx_st3_hvalid
		output wire          pio_tx_st3_pvalid_o       //                 .tx_st3_pvalid
	);

	intel_pcie_bam_v2_hwtcl #(
		.VFNUM_WIDTH   (12),
		.PFNUM_WIDTH   (2),
		.DATA_WIDTH    (1024),
		.DEVICE_FAMILY ("Agilex")
	) pio0 (
		.Clk_i                    (Clk_i),                    //   input,     width = 1,              clk.clk
		.Rstn_i                   (Rstn_i),                   //   input,     width = 1,            reset.reset_n
		.pio_clk                  (pio_clk),                  //  output,     width = 1,   pio_master_clk.clk
		.pio_rst_n                (pio_rst_n),                //  output,     width = 1, pio_master_reset.reset_n
		.pio_address_o            (pio_address_o),            //  output,    width = 64,       pio_master.address
		.pio_read_o               (pio_read_o),               //  output,     width = 1,                 .read
		.pio_readdata_i           (pio_readdata_i),           //   input,  width = 1024,                 .readdata
		.pio_readdatavalid_i      (pio_readdatavalid_i),      //   input,     width = 1,                 .readdatavalid
		.pio_write_o              (pio_write_o),              //  output,     width = 1,                 .write
		.pio_writedata_o          (pio_writedata_o),          //  output,  width = 1024,                 .writedata
		.pio_waitrequest_i        (pio_waitrequest_i),        //   input,     width = 1,                 .waitrequest
		.pio_byteenable_o         (pio_byteenable_o),         //  output,   width = 128,                 .byteenable
		.pio_response_i           (pio_response_i),           //   input,     width = 2,                 .response
		.pio_burstcount_o         (pio_burstcount_o),         //  output,     width = 4,                 .burstcount
		.pio_rx_st0_payload_i     (pio_rx_st0_payload_i),     //   input,   width = 256,       rx_st0_pio.data
		.pio_rx_st0_sop_i         (pio_rx_st0_sop_i),         //   input,     width = 1,                 .startofpacket
		.pio_rx_st0_eop_i         (pio_rx_st0_eop_i),         //   input,     width = 1,                 .endofpacket
		.pio_rx_st0_dvalid_i      (pio_rx_st0_dvalid_i),      //   input,     width = 1,                 .valid
		.pio_rx_st0_empty_i       (pio_rx_st0_empty_i),       //   input,     width = 3,                 .empty
		.pio_rx_st_ready_o        (pio_rx_st_ready_o),        //  output,     width = 1,                 .ready
		.pio_rx_st1_payload_i     (pio_rx_st1_payload_i),     //   input,   width = 256,       rx_st1_pio.data
		.pio_rx_st1_sop_i         (pio_rx_st1_sop_i),         //   input,     width = 1,                 .startofpacket
		.pio_rx_st1_eop_i         (pio_rx_st1_eop_i),         //   input,     width = 1,                 .endofpacket
		.pio_rx_st1_dvalid_i      (pio_rx_st1_dvalid_i),      //   input,     width = 1,                 .valid
		.pio_rx_st1_empty_i       (pio_rx_st1_empty_i),       //   input,     width = 3,                 .empty
		.pio_rx_st2_payload_i     (pio_rx_st2_payload_i),     //   input,   width = 256,       rx_st2_pio.data
		.pio_rx_st2_sop_i         (pio_rx_st2_sop_i),         //   input,     width = 1,                 .startofpacket
		.pio_rx_st2_eop_i         (pio_rx_st2_eop_i),         //   input,     width = 1,                 .endofpacket
		.pio_rx_st2_dvalid_i      (pio_rx_st2_dvalid_i),      //   input,     width = 1,                 .valid
		.pio_rx_st2_empty_i       (pio_rx_st2_empty_i),       //   input,     width = 3,                 .empty
		.pio_rx_st3_payload_i     (pio_rx_st3_payload_i),     //   input,   width = 256,       rx_st3_pio.data
		.pio_rx_st3_sop_i         (pio_rx_st3_sop_i),         //   input,     width = 1,                 .startofpacket
		.pio_rx_st3_eop_i         (pio_rx_st3_eop_i),         //   input,     width = 1,                 .endofpacket
		.pio_rx_st3_dvalid_i      (pio_rx_st3_dvalid_i),      //   input,     width = 1,                 .valid
		.pio_rx_st3_empty_i       (pio_rx_st3_empty_i),       //   input,     width = 3,                 .empty
		.rx_st_hcrdt_init_o       (rx_st_hcrdt_init_o),       //  output,     width = 3,  rx_st0_pio_misc.rx_st_Hcrdt_init
		.rx_st_hcrdt_update_o     (rx_st_hcrdt_update_o),     //  output,     width = 3,                 .rx_st_Hcrdt_update
		.rx_st_hcrdt_update_cnt_o (rx_st_hcrdt_update_cnt_o), //  output,     width = 6,                 .rx_st_Hcrdt_update_cnt
		.rx_st_hcrdt_init_ack_i   (rx_st_hcrdt_init_ack_i),   //   input,     width = 3,                 .rx_st_Hcrdt_init_ack
		.rx_st_dcrdt_init_o       (rx_st_dcrdt_init_o),       //  output,     width = 3,                 .rx_st_Dcrdt_init
		.rx_st_dcrdt_update_o     (rx_st_dcrdt_update_o),     //  output,     width = 3,                 .rx_st_Dcrdt_update
		.rx_st_dcrdt_update_cnt_o (rx_st_dcrdt_update_cnt_o), //  output,    width = 12,                 .rx_st_Dcrdt_update_cnt
		.rx_st_dcrdt_init_ack_i   (rx_st_dcrdt_init_ack_i),   //   input,     width = 3,                 .rx_st_Dcrdt_init_ack
		.pio_rx_st0_header_i      (pio_rx_st0_header_i),      //   input,   width = 128,                 .rx_st0_hdr
		.pio_rx_st0_tlp_prfx_i    (pio_rx_st0_tlp_prfx_i),    //   input,    width = 32,                 .rx_st0_prefix
		.pio_rx_st0_hvalid_i      (pio_rx_st0_hvalid_i),      //   input,     width = 1,                 .rx_st0_hvalid
		.pio_rx_st0_pvalid_i      (pio_rx_st0_pvalid_i),      //   input,     width = 1,                 .rx_st0_pvalid
		.pio_rx_st0_bar_i         (pio_rx_st0_bar_i),         //   input,     width = 3,                 .rx_st0_bar
		.pio_rx_st1_header_i      (pio_rx_st1_header_i),      //   input,   width = 128,                 .rx_st1_hdr
		.pio_rx_st1_tlp_prfx_i    (pio_rx_st1_tlp_prfx_i),    //   input,    width = 32,                 .rx_st1_prefix
		.pio_rx_st1_hvalid_i      (pio_rx_st1_hvalid_i),      //   input,     width = 1,                 .rx_st1_hvalid
		.pio_rx_st1_pvalid_i      (pio_rx_st1_pvalid_i),      //   input,     width = 1,                 .rx_st1_pvalid
		.pio_rx_st1_bar_i         (pio_rx_st1_bar_i),         //   input,     width = 3,                 .rx_st1_bar
		.pio_rx_st2_header_i      (pio_rx_st2_header_i),      //   input,   width = 128,                 .rx_st2_hdr
		.pio_rx_st2_tlp_prfx_i    (pio_rx_st2_tlp_prfx_i),    //   input,    width = 32,                 .rx_st2_prefix
		.pio_rx_st2_hvalid_i      (pio_rx_st2_hvalid_i),      //   input,     width = 1,                 .rx_st2_hvalid
		.pio_rx_st2_pvalid_i      (pio_rx_st2_pvalid_i),      //   input,     width = 1,                 .rx_st2_pvalid
		.pio_rx_st2_bar_i         (pio_rx_st2_bar_i),         //   input,     width = 3,                 .rx_st2_bar
		.pio_rx_st3_header_i      (pio_rx_st3_header_i),      //   input,   width = 128,                 .rx_st3_hdr
		.pio_rx_st3_tlp_prfx_i    (pio_rx_st3_tlp_prfx_i),    //   input,    width = 32,                 .rx_st3_prefix
		.pio_rx_st3_hvalid_i      (pio_rx_st3_hvalid_i),      //   input,     width = 1,                 .rx_st3_hvalid
		.pio_rx_st3_pvalid_i      (pio_rx_st3_pvalid_i),      //   input,     width = 1,                 .rx_st3_pvalid
		.pio_rx_st3_bar_i         (pio_rx_st3_bar_i),         //   input,     width = 3,                 .rx_st3_bar
		.pio_tx_st0_payload_o     (pio_tx_st0_payload_o),     //  output,   width = 256,       tx_st0_pio.data
		.pio_tx_st0_sop_o         (pio_tx_st0_sop_o),         //  output,     width = 1,                 .startofpacket
		.pio_tx_st0_eop_o         (pio_tx_st0_eop_o),         //  output,     width = 1,                 .endofpacket
		.pio_tx_st0_dvalid_o      (pio_tx_st0_dvalid_o),      //  output,     width = 1,                 .valid
		.pio_tx_st_ready_i        (pio_tx_st_ready_i),        //   input,     width = 1,                 .ready
		.pio_tx_st1_payload_o     (pio_tx_st1_payload_o),     //  output,   width = 256,       tx_st1_pio.data
		.pio_tx_st1_sop_o         (pio_tx_st1_sop_o),         //  output,     width = 1,                 .startofpacket
		.pio_tx_st1_eop_o         (pio_tx_st1_eop_o),         //  output,     width = 1,                 .endofpacket
		.pio_tx_st1_dvalid_o      (pio_tx_st1_dvalid_o),      //  output,     width = 1,                 .valid
		.pio_tx_st2_payload_o     (pio_tx_st2_payload_o),     //  output,   width = 256,       tx_st2_pio.data
		.pio_tx_st2_sop_o         (pio_tx_st2_sop_o),         //  output,     width = 1,                 .startofpacket
		.pio_tx_st2_eop_o         (pio_tx_st2_eop_o),         //  output,     width = 1,                 .endofpacket
		.pio_tx_st2_dvalid_o      (pio_tx_st2_dvalid_o),      //  output,     width = 1,                 .valid
		.pio_tx_st3_payload_o     (pio_tx_st3_payload_o),     //  output,   width = 256,       tx_st3_pio.data
		.pio_tx_st3_sop_o         (pio_tx_st3_sop_o),         //  output,     width = 1,                 .startofpacket
		.pio_tx_st3_eop_o         (pio_tx_st3_eop_o),         //  output,     width = 1,                 .endofpacket
		.pio_tx_st3_dvalid_o      (pio_tx_st3_dvalid_o),      //  output,     width = 1,                 .valid
		.pio_tx_st0_header_o      (pio_tx_st0_header_o),      //  output,   width = 128,  tx_st0_pio_misc.tx_st0_hdr
		.pio_tx_st1_header_o      (pio_tx_st1_header_o),      //  output,   width = 128,                 .tx_st1_hdr
		.pio_tx_st2_header_o      (pio_tx_st2_header_o),      //  output,   width = 128,                 .tx_st2_hdr
		.pio_tx_st3_header_o      (pio_tx_st3_header_o),      //  output,   width = 128,                 .tx_st3_hdr
		.tx_st_hcrdt_init_i       (tx_st_hcrdt_init_i),       //   input,     width = 3,                 .tx_st_Hcrdt_init
		.tx_st_hcrdt_update_i     (tx_st_hcrdt_update_i),     //   input,     width = 3,                 .tx_st_Hcrdt_update
		.tx_st_hcrdt_update_cnt_i (tx_st_hcrdt_update_cnt_i), //   input,     width = 6,                 .tx_st_Hcrdt_update_cnt
		.tx_st_hcrdt_init_ack_o   (tx_st_hcrdt_init_ack_o),   //  output,     width = 3,                 .tx_st_Hcrdtt_init_ack
		.tx_st_dcrdt_init_i       (tx_st_dcrdt_init_i),       //   input,     width = 3,                 .tx_st_Dcrdt_init
		.tx_st_dcrdt_update_i     (tx_st_dcrdt_update_i),     //   input,     width = 3,                 .tx_st_Dcrdt_update
		.tx_st_dcrdt_update_cnt_i (tx_st_dcrdt_update_cnt_i), //   input,    width = 12,                 .tx_st_Dcrdt_update_cnt
		.tx_st_dcrdt_init_ack_o   (tx_st_dcrdt_init_ack_o),   //  output,     width = 3,                 .tx_st_Dcrdt_init_ack
		.pio_tx_st0_prefix_o      (pio_tx_st0_prefix_o),      //  output,    width = 32,                 .tx_st0_prefix
		.pio_tx_st0_hvalid_o      (pio_tx_st0_hvalid_o),      //  output,     width = 1,                 .tx_st0_hvalid
		.pio_tx_st0_pvalid_o      (pio_tx_st0_pvalid_o),      //  output,     width = 1,                 .tx_st0_pvalid
		.pio_tx_st1_prefix_o      (pio_tx_st1_prefix_o),      //  output,    width = 32,                 .tx_st1_prefix
		.pio_tx_st1_hvalid_o      (pio_tx_st1_hvalid_o),      //  output,     width = 1,                 .tx_st1_hvalid
		.pio_tx_st1_pvalid_o      (pio_tx_st1_pvalid_o),      //  output,     width = 1,                 .tx_st1_pvalid
		.pio_tx_st2_prefix_o      (pio_tx_st2_prefix_o),      //  output,    width = 32,                 .tx_st2_prefix
		.pio_tx_st2_hvalid_o      (pio_tx_st2_hvalid_o),      //  output,     width = 1,                 .tx_st2_hvalid
		.pio_tx_st2_pvalid_o      (pio_tx_st2_pvalid_o),      //  output,     width = 1,                 .tx_st2_pvalid
		.pio_tx_st3_prefix_o      (pio_tx_st3_prefix_o),      //  output,    width = 32,                 .tx_st3_prefix
		.pio_tx_st3_hvalid_o      (pio_tx_st3_hvalid_o),      //  output,     width = 1,                 .tx_st3_hvalid
		.pio_tx_st3_pvalid_o      (pio_tx_st3_pvalid_o)       //  output,     width = 1,                 .tx_st3_pvalid
	);

endmodule
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "EtAh8aN7m2BPKOTfO5tEAbNSD19BnNEklF4xQRY7YZ2oRe/8wDIRx8XCKuwkXQtjYcM5gRXSD6c+oGX77mfnvlAGw9KTmnXPBu3GU7e3qFjUTrXWlEAN76gMqJTePk91Iv2qtpAKuY2LJHLiowUVDoSuAt1Csh1O2u7qDzQRIaeVL/AJWYDMfWERE2K26wZcHHB8eTbMnhSND4m01aQODfKXixyUFYBUVJCy/gZrUwDeZiH4XE6JthCMbIphHj+XrJk6umYqQBuFOenzn2gOMXR7PeNe89DBDQ4hTBT+o43WAVV4QxqLIdiXcMS2px5DRDRHf8N2b2HEoBv+zuCeyXjSRAUXxw+N4o2BGpUSLr0oM3Omm9pjwYGrUd5sVRe3jFY9zU4jAcB2BZu29c2viQwJlHJqyYed0vLXCPFZb1ODr5wYL4wJOZgcuTk4jcEmZvGktMaJDL8xCH4UA5ymUVpXy3eT7Oh+jlASkcAwK55LyjlOUjH6mt9ssfG1oEUpN/zG8JMu+UTp8h9T7ZKyNlbY0UKwXthkYQ7BNM8xH0JhawWxonq5ed23j8zVe8XVH7QXH4nVodl56W0VeJ0qbZa8JsTZK1a0MkGFS2peDOyIDIEfaBPAnfsuvni6IygXA9SrNmpNJKyG2sDqNaNyBQV9hdgm/q+BueW/0vR207hDNQ+VIBuIbMRJo8YgBMINOva08gRnOXV9jScE/Ai9Qo2YaMijcq0EMG64VrltjN1vBHs6FAWxKrhYZ/ge1LJikyQKWV14mIHlhGwcgB6WoTb5WJuFJfShXlInh/31bZnOJpPi2tYqthpnEaVe+7Ub5kDPOpS5v2FPMidFkb5/H5G1MjL8ib32YIR+MV/NvkgE0+yISBW216GWj23y68SsZ4iXdpGcLgwrVZI92X8a9k4IbrX8bGo6A5FrnpSwmZN1RFD5kOE0aPC34yvLhNKdhj+zBChDpD4wpZP2Z9N403N+7TYBKeILm2XZLvVHaIVM9/HWVCZhCANcIfqNB/XZ"
`endif