// (C) 2001-2023 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


// Copyright 2022 Intel Corporation.
//
// THIS SOFTWARE MAY CONTAIN PREPRODUCTION CODE AND IS PROVIDED BY THE
// COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS OR IMPLIED
// WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF
// MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE
// LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
// SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR
// BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY,
// WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE
// OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE,
// EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
///////////////////////////////////////////////////////////////////////

//-------------------------------------------------------------------------
//  Global Defines
// ------------------------------------------------------------------------
//

`ifndef CXLTYP2_DEFINES
`define CXLTYP2_DEFINES


package cxl_type2_defines;



    //# HDL Defines
    //# =====================

    `define LVF2
    `define QUARTUS_FPGA_SYNTH
    `define INCLUDE_CXLMEM_READY //?
    `define ENABLE_DDR_DBI_PINS //?
    `define HDM_16G 
    `define SPR_D0
    `define SUPPORT_ALGORITHM_1A
    `define ALG_1A_SUPPORT_SELF_CHECK
    `define RNR_B0_TILE 
    `define ENABLE_1_BBS_SLICE


   `define OOO_SUPPORT
   `define OOORSP
   `define OOORSP_MC_AXI2AVMM

// For user reference:
// `ifdef SPR_A0
//  assign POR_BBS_DCCCFG.SPRBUG_m2smetafield  = 1'b1;
//  assign POR_BBS_DCCCFG.SPRBUG_m2smeminvcmpe = 1'b1;
//  assign POR_BBS_DCCCFG.SPRBUG_m2swrsnpinva  = 1'b0;
//`elsif SPR_B0
//  assign POR_BBS_DCCCFG.SPRBUG_m2smetafield  = 1'b0;
//  assign POR_BBS_DCCCFG.SPRBUG_m2smeminvcmpe = 1'b1;
//  assign POR_BBS_DCCCFG.SPRBUG_m2swrsnpinva  = 1'b0;
//`elsif SPR_D0
//  assign POR_BBS_DCCCFG.SPRBUG_m2smetafield  = 1'b0;
//  assign POR_BBS_DCCCFG.SPRBUG_m2smeminvcmpe = 1'b0;
//  assign POR_BBS_DCCCFG.SPRBUG_m2swrsnpinva  = 1'b1;
//`else
//  assign POR_BBS_DCCCFG.SPRBUG_m2smetafield  = 1'b0;
//  assign POR_BBS_DCCCFG.SPRBUG_m2smeminvcmpe = 1'b0;
//  assign POR_BBS_DCCCFG.SPRBUG_m2swrsnpinva  = 1'b0;
//`endif

endpackage
`endif// `define CXLTYP2_DEFINES

