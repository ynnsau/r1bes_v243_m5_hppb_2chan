// (C) 2001-2024 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


// pcie_ed_altera_mm_interconnect_1920_sx2feoa.v

// This file was auto-generated from altera_mm_interconnect_hw.tcl.  If you edit it your changes
// will probably be lost.
// 
// Generated using ACDS version 22.1 174

`timescale 1 ps / 1 ps
module pcie_ed_altera_mm_interconnect_1920_sx2feoa (
		input  wire [63:0]   pio0_pio_master_address,                                      //                                        pio0_pio_master.address
		output wire          pio0_pio_master_waitrequest,                                  //                                                       .waitrequest
		input  wire [3:0]    pio0_pio_master_burstcount,                                   //                                                       .burstcount
		input  wire [127:0]  pio0_pio_master_byteenable,                                   //                                                       .byteenable
		input  wire          pio0_pio_master_read,                                         //                                                       .read
		output wire [1023:0] pio0_pio_master_readdata,                                     //                                                       .readdata
		output wire          pio0_pio_master_readdatavalid,                                //                                                       .readdatavalid
		input  wire          pio0_pio_master_write,                                        //                                                       .write
		input  wire [1023:0] pio0_pio_master_writedata,                                    //                                                       .writedata
		output wire [1:0]    pio0_pio_master_response,                                     //                                                       .response
		output wire [7:0]    MEM0_s1_address,                                              //                                                MEM0_s1.address
		output wire          MEM0_s1_write,                                                //                                                       .write
		input  wire [1023:0] MEM0_s1_readdata,                                             //                                                       .readdata
		output wire [1023:0] MEM0_s1_writedata,                                            //                                                       .writedata
		output wire [127:0]  MEM0_s1_byteenable,                                           //                                                       .byteenable
		output wire          MEM0_s1_chipselect,                                           //                                                       .chipselect
		output wire          MEM0_s1_clken,                                                //                                                       .clken
		input  wire          MEM0_reset1_reset_bridge_in_reset_reset,                      //                      MEM0_reset1_reset_bridge_in_reset.reset
		input  wire          pio0_pio_master_translator_reset_reset_bridge_in_reset_reset, // pio0_pio_master_translator_reset_reset_bridge_in_reset.reset
		input  wire          pio0_pio_master_clk_clk                                       //                                    pio0_pio_master_clk.clk
	);

	wire           pio0_pio_master_translator_avalon_universal_master_0_waitrequest;   // pio0_pio_master_agent:av_waitrequest -> pio0_pio_master_translator:uav_waitrequest
	wire  [1023:0] pio0_pio_master_translator_avalon_universal_master_0_readdata;      // pio0_pio_master_agent:av_readdata -> pio0_pio_master_translator:uav_readdata
	wire           pio0_pio_master_translator_avalon_universal_master_0_debugaccess;   // pio0_pio_master_translator:uav_debugaccess -> pio0_pio_master_agent:av_debugaccess
	wire    [63:0] pio0_pio_master_translator_avalon_universal_master_0_address;       // pio0_pio_master_translator:uav_address -> pio0_pio_master_agent:av_address
	wire           pio0_pio_master_translator_avalon_universal_master_0_read;          // pio0_pio_master_translator:uav_read -> pio0_pio_master_agent:av_read
	wire   [127:0] pio0_pio_master_translator_avalon_universal_master_0_byteenable;    // pio0_pio_master_translator:uav_byteenable -> pio0_pio_master_agent:av_byteenable
	wire           pio0_pio_master_translator_avalon_universal_master_0_readdatavalid; // pio0_pio_master_agent:av_readdatavalid -> pio0_pio_master_translator:uav_readdatavalid
	wire     [1:0] pio0_pio_master_translator_avalon_universal_master_0_response;      // pio0_pio_master_agent:av_response -> pio0_pio_master_translator:uav_response
	wire           pio0_pio_master_translator_avalon_universal_master_0_lock;          // pio0_pio_master_translator:uav_lock -> pio0_pio_master_agent:av_lock
	wire           pio0_pio_master_translator_avalon_universal_master_0_write;         // pio0_pio_master_translator:uav_write -> pio0_pio_master_agent:av_write
	wire  [1023:0] pio0_pio_master_translator_avalon_universal_master_0_writedata;     // pio0_pio_master_translator:uav_writedata -> pio0_pio_master_agent:av_writedata
	wire    [10:0] pio0_pio_master_translator_avalon_universal_master_0_burstcount;    // pio0_pio_master_translator:uav_burstcount -> pio0_pio_master_agent:av_burstcount
	wire           rsp_mux_src_valid;                                                  // rsp_mux:src_valid -> pio0_pio_master_agent:rp_valid
	wire  [1266:0] rsp_mux_src_data;                                                   // rsp_mux:src_data -> pio0_pio_master_agent:rp_data
	wire           rsp_mux_src_ready;                                                  // pio0_pio_master_agent:rp_ready -> rsp_mux:src_ready
	wire     [0:0] rsp_mux_src_channel;                                                // rsp_mux:src_channel -> pio0_pio_master_agent:rp_channel
	wire           rsp_mux_src_startofpacket;                                          // rsp_mux:src_startofpacket -> pio0_pio_master_agent:rp_startofpacket
	wire           rsp_mux_src_endofpacket;                                            // rsp_mux:src_endofpacket -> pio0_pio_master_agent:rp_endofpacket
	wire  [1023:0] mem0_s1_agent_m0_readdata;                                          // MEM0_s1_translator:uav_readdata -> MEM0_s1_agent:m0_readdata
	wire           mem0_s1_agent_m0_waitrequest;                                       // MEM0_s1_translator:uav_waitrequest -> MEM0_s1_agent:m0_waitrequest
	wire           mem0_s1_agent_m0_debugaccess;                                       // MEM0_s1_agent:m0_debugaccess -> MEM0_s1_translator:uav_debugaccess
	wire    [63:0] mem0_s1_agent_m0_address;                                           // MEM0_s1_agent:m0_address -> MEM0_s1_translator:uav_address
	wire   [127:0] mem0_s1_agent_m0_byteenable;                                        // MEM0_s1_agent:m0_byteenable -> MEM0_s1_translator:uav_byteenable
	wire           mem0_s1_agent_m0_read;                                              // MEM0_s1_agent:m0_read -> MEM0_s1_translator:uav_read
	wire           mem0_s1_agent_m0_readdatavalid;                                     // MEM0_s1_translator:uav_readdatavalid -> MEM0_s1_agent:m0_readdatavalid
	wire           mem0_s1_agent_m0_lock;                                              // MEM0_s1_agent:m0_lock -> MEM0_s1_translator:uav_lock
	wire  [1023:0] mem0_s1_agent_m0_writedata;                                         // MEM0_s1_agent:m0_writedata -> MEM0_s1_translator:uav_writedata
	wire           mem0_s1_agent_m0_write;                                             // MEM0_s1_agent:m0_write -> MEM0_s1_translator:uav_write
	wire     [7:0] mem0_s1_agent_m0_burstcount;                                        // MEM0_s1_agent:m0_burstcount -> MEM0_s1_translator:uav_burstcount
	wire           mem0_s1_agent_rf_source_valid;                                      // MEM0_s1_agent:rf_source_valid -> MEM0_s1_agent_rsp_fifo:in_valid
	wire  [1267:0] mem0_s1_agent_rf_source_data;                                       // MEM0_s1_agent:rf_source_data -> MEM0_s1_agent_rsp_fifo:in_data
	wire           mem0_s1_agent_rf_source_ready;                                      // MEM0_s1_agent_rsp_fifo:in_ready -> MEM0_s1_agent:rf_source_ready
	wire           mem0_s1_agent_rf_source_startofpacket;                              // MEM0_s1_agent:rf_source_startofpacket -> MEM0_s1_agent_rsp_fifo:in_startofpacket
	wire           mem0_s1_agent_rf_source_endofpacket;                                // MEM0_s1_agent:rf_source_endofpacket -> MEM0_s1_agent_rsp_fifo:in_endofpacket
	wire           mem0_s1_agent_rsp_fifo_out_valid;                                   // MEM0_s1_agent_rsp_fifo:out_valid -> MEM0_s1_agent:rf_sink_valid
	wire  [1267:0] mem0_s1_agent_rsp_fifo_out_data;                                    // MEM0_s1_agent_rsp_fifo:out_data -> MEM0_s1_agent:rf_sink_data
	wire           mem0_s1_agent_rsp_fifo_out_ready;                                   // MEM0_s1_agent:rf_sink_ready -> MEM0_s1_agent_rsp_fifo:out_ready
	wire           mem0_s1_agent_rsp_fifo_out_startofpacket;                           // MEM0_s1_agent_rsp_fifo:out_startofpacket -> MEM0_s1_agent:rf_sink_startofpacket
	wire           mem0_s1_agent_rsp_fifo_out_endofpacket;                             // MEM0_s1_agent_rsp_fifo:out_endofpacket -> MEM0_s1_agent:rf_sink_endofpacket
	wire           mem0_s1_agent_rdata_fifo_src_valid;                                 // MEM0_s1_agent:rdata_fifo_src_valid -> MEM0_s1_agent:rdata_fifo_sink_valid
	wire  [1025:0] mem0_s1_agent_rdata_fifo_src_data;                                  // MEM0_s1_agent:rdata_fifo_src_data -> MEM0_s1_agent:rdata_fifo_sink_data
	wire           mem0_s1_agent_rdata_fifo_src_ready;                                 // MEM0_s1_agent:rdata_fifo_sink_ready -> MEM0_s1_agent:rdata_fifo_src_ready
	wire           pio0_pio_master_agent_cp_valid;                                     // pio0_pio_master_agent:cp_valid -> router:sink_valid
	wire  [1266:0] pio0_pio_master_agent_cp_data;                                      // pio0_pio_master_agent:cp_data -> router:sink_data
	wire           pio0_pio_master_agent_cp_ready;                                     // router:sink_ready -> pio0_pio_master_agent:cp_ready
	wire           pio0_pio_master_agent_cp_startofpacket;                             // pio0_pio_master_agent:cp_startofpacket -> router:sink_startofpacket
	wire           pio0_pio_master_agent_cp_endofpacket;                               // pio0_pio_master_agent:cp_endofpacket -> router:sink_endofpacket
	wire           router_src_valid;                                                   // router:src_valid -> cmd_demux:sink_valid
	wire  [1266:0] router_src_data;                                                    // router:src_data -> cmd_demux:sink_data
	wire           router_src_ready;                                                   // cmd_demux:sink_ready -> router:src_ready
	wire     [0:0] router_src_channel;                                                 // router:src_channel -> cmd_demux:sink_channel
	wire           router_src_startofpacket;                                           // router:src_startofpacket -> cmd_demux:sink_startofpacket
	wire           router_src_endofpacket;                                             // router:src_endofpacket -> cmd_demux:sink_endofpacket
	wire           mem0_s1_agent_rp_valid;                                             // MEM0_s1_agent:rp_valid -> router_001:sink_valid
	wire  [1266:0] mem0_s1_agent_rp_data;                                              // MEM0_s1_agent:rp_data -> router_001:sink_data
	wire           mem0_s1_agent_rp_ready;                                             // router_001:sink_ready -> MEM0_s1_agent:rp_ready
	wire           mem0_s1_agent_rp_startofpacket;                                     // MEM0_s1_agent:rp_startofpacket -> router_001:sink_startofpacket
	wire           mem0_s1_agent_rp_endofpacket;                                       // MEM0_s1_agent:rp_endofpacket -> router_001:sink_endofpacket
	wire           router_001_src_valid;                                               // router_001:src_valid -> rsp_demux:sink_valid
	wire  [1266:0] router_001_src_data;                                                // router_001:src_data -> rsp_demux:sink_data
	wire           router_001_src_ready;                                               // rsp_demux:sink_ready -> router_001:src_ready
	wire     [0:0] router_001_src_channel;                                             // router_001:src_channel -> rsp_demux:sink_channel
	wire           router_001_src_startofpacket;                                       // router_001:src_startofpacket -> rsp_demux:sink_startofpacket
	wire           router_001_src_endofpacket;                                         // router_001:src_endofpacket -> rsp_demux:sink_endofpacket
	wire           cmd_mux_src_valid;                                                  // cmd_mux:src_valid -> MEM0_s1_burst_adapter:sink0_valid
	wire  [1266:0] cmd_mux_src_data;                                                   // cmd_mux:src_data -> MEM0_s1_burst_adapter:sink0_data
	wire           cmd_mux_src_ready;                                                  // MEM0_s1_burst_adapter:sink0_ready -> cmd_mux:src_ready
	wire     [0:0] cmd_mux_src_channel;                                                // cmd_mux:src_channel -> MEM0_s1_burst_adapter:sink0_channel
	wire           cmd_mux_src_startofpacket;                                          // cmd_mux:src_startofpacket -> MEM0_s1_burst_adapter:sink0_startofpacket
	wire           cmd_mux_src_endofpacket;                                            // cmd_mux:src_endofpacket -> MEM0_s1_burst_adapter:sink0_endofpacket
	wire           mem0_s1_burst_adapter_source0_valid;                                // MEM0_s1_burst_adapter:source0_valid -> MEM0_s1_agent:cp_valid
	wire  [1266:0] mem0_s1_burst_adapter_source0_data;                                 // MEM0_s1_burst_adapter:source0_data -> MEM0_s1_agent:cp_data
	wire           mem0_s1_burst_adapter_source0_ready;                                // MEM0_s1_agent:cp_ready -> MEM0_s1_burst_adapter:source0_ready
	wire     [0:0] mem0_s1_burst_adapter_source0_channel;                              // MEM0_s1_burst_adapter:source0_channel -> MEM0_s1_agent:cp_channel
	wire           mem0_s1_burst_adapter_source0_startofpacket;                        // MEM0_s1_burst_adapter:source0_startofpacket -> MEM0_s1_agent:cp_startofpacket
	wire           mem0_s1_burst_adapter_source0_endofpacket;                          // MEM0_s1_burst_adapter:source0_endofpacket -> MEM0_s1_agent:cp_endofpacket
	wire           cmd_demux_src0_valid;                                               // cmd_demux:src0_valid -> cmd_mux:sink0_valid
	wire  [1266:0] cmd_demux_src0_data;                                                // cmd_demux:src0_data -> cmd_mux:sink0_data
	wire           cmd_demux_src0_ready;                                               // cmd_mux:sink0_ready -> cmd_demux:src0_ready
	wire     [0:0] cmd_demux_src0_channel;                                             // cmd_demux:src0_channel -> cmd_mux:sink0_channel
	wire           cmd_demux_src0_startofpacket;                                       // cmd_demux:src0_startofpacket -> cmd_mux:sink0_startofpacket
	wire           cmd_demux_src0_endofpacket;                                         // cmd_demux:src0_endofpacket -> cmd_mux:sink0_endofpacket
	wire           rsp_demux_src0_valid;                                               // rsp_demux:src0_valid -> rsp_mux:sink0_valid
	wire  [1266:0] rsp_demux_src0_data;                                                // rsp_demux:src0_data -> rsp_mux:sink0_data
	wire           rsp_demux_src0_ready;                                               // rsp_mux:sink0_ready -> rsp_demux:src0_ready
	wire     [0:0] rsp_demux_src0_channel;                                             // rsp_demux:src0_channel -> rsp_mux:sink0_channel
	wire           rsp_demux_src0_startofpacket;                                       // rsp_demux:src0_startofpacket -> rsp_mux:sink0_startofpacket
	wire           rsp_demux_src0_endofpacket;                                         // rsp_demux:src0_endofpacket -> rsp_mux:sink0_endofpacket

	pcie_ed_altera_merlin_master_translator_191_g7h47bq #(
		.AV_ADDRESS_W                (64),
		.AV_DATA_W                   (1024),
		.AV_BURSTCOUNT_W             (4),
		.AV_BYTEENABLE_W             (128),
		.UAV_ADDRESS_W               (64),
		.UAV_BURSTCOUNT_W            (11),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (1),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (128),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (1),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0),
		.SYNC_RESET                  (1),
		.WAITREQUEST_ALLOWANCE       (0)
	) pio0_pio_master_translator (
		.clk                    (pio0_pio_master_clk_clk),                                            //   input,     width = 1,                       clk.clk
		.reset                  (pio0_pio_master_translator_reset_reset_bridge_in_reset_reset),       //   input,     width = 1,                     reset.reset
		.uav_address            (pio0_pio_master_translator_avalon_universal_master_0_address),       //  output,    width = 64, avalon_universal_master_0.address
		.uav_burstcount         (pio0_pio_master_translator_avalon_universal_master_0_burstcount),    //  output,    width = 11,                          .burstcount
		.uav_read               (pio0_pio_master_translator_avalon_universal_master_0_read),          //  output,     width = 1,                          .read
		.uav_write              (pio0_pio_master_translator_avalon_universal_master_0_write),         //  output,     width = 1,                          .write
		.uav_waitrequest        (pio0_pio_master_translator_avalon_universal_master_0_waitrequest),   //   input,     width = 1,                          .waitrequest
		.uav_readdatavalid      (pio0_pio_master_translator_avalon_universal_master_0_readdatavalid), //   input,     width = 1,                          .readdatavalid
		.uav_byteenable         (pio0_pio_master_translator_avalon_universal_master_0_byteenable),    //  output,   width = 128,                          .byteenable
		.uav_readdata           (pio0_pio_master_translator_avalon_universal_master_0_readdata),      //   input,  width = 1024,                          .readdata
		.uav_writedata          (pio0_pio_master_translator_avalon_universal_master_0_writedata),     //  output,  width = 1024,                          .writedata
		.uav_lock               (pio0_pio_master_translator_avalon_universal_master_0_lock),          //  output,     width = 1,                          .lock
		.uav_debugaccess        (pio0_pio_master_translator_avalon_universal_master_0_debugaccess),   //  output,     width = 1,                          .debugaccess
		.uav_response           (pio0_pio_master_translator_avalon_universal_master_0_response),      //   input,     width = 2,                          .response
		.av_address             (pio0_pio_master_address),                                            //   input,    width = 64,      avalon_anti_master_0.address
		.av_waitrequest         (pio0_pio_master_waitrequest),                                        //  output,     width = 1,                          .waitrequest
		.av_burstcount          (pio0_pio_master_burstcount),                                         //   input,     width = 4,                          .burstcount
		.av_byteenable          (pio0_pio_master_byteenable),                                         //   input,   width = 128,                          .byteenable
		.av_read                (pio0_pio_master_read),                                               //   input,     width = 1,                          .read
		.av_readdata            (pio0_pio_master_readdata),                                           //  output,  width = 1024,                          .readdata
		.av_readdatavalid       (pio0_pio_master_readdatavalid),                                      //  output,     width = 1,                          .readdatavalid
		.av_write               (pio0_pio_master_write),                                              //   input,     width = 1,                          .write
		.av_writedata           (pio0_pio_master_writedata),                                          //   input,  width = 1024,                          .writedata
		.av_response            (pio0_pio_master_response),                                           //  output,     width = 2,                          .response
		.av_beginbursttransfer  (1'b0),                                                               // (terminated),                                          
		.av_begintransfer       (1'b0),                                                               // (terminated),                                          
		.av_chipselect          (1'b0),                                                               // (terminated),                                          
		.av_lock                (1'b0),                                                               // (terminated),                                          
		.av_debugaccess         (1'b0),                                                               // (terminated),                                          
		.uav_clken              (),                                                                   // (terminated),                                          
		.av_clken               (1'b1),                                                               // (terminated),                                          
		.uav_writeresponsevalid (1'b0),                                                               // (terminated),                                          
		.av_writeresponsevalid  ()                                                                    // (terminated),                                          
	);

	pcie_ed_altera_merlin_slave_translator_191_x56fcki #(
		.AV_ADDRESS_W                   (8),
		.AV_DATA_W                      (1024),
		.UAV_DATA_W                     (1024),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (128),
		.UAV_BYTEENABLE_W               (128),
		.UAV_ADDRESS_W                  (64),
		.UAV_BURSTCOUNT_W               (8),
		.AV_READLATENCY                 (2),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (128),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0),
		.WAITREQUEST_ALLOWANCE          (0),
		.SYNC_RESET                     (1)
	) mem0_s1_translator (
		.clk                    (pio0_pio_master_clk_clk),                                      //   input,     width = 1,                      clk.clk
		.reset                  (pio0_pio_master_translator_reset_reset_bridge_in_reset_reset), //   input,     width = 1,                    reset.reset
		.uav_address            (mem0_s1_agent_m0_address),                                     //   input,    width = 64, avalon_universal_slave_0.address
		.uav_burstcount         (mem0_s1_agent_m0_burstcount),                                  //   input,     width = 8,                         .burstcount
		.uav_read               (mem0_s1_agent_m0_read),                                        //   input,     width = 1,                         .read
		.uav_write              (mem0_s1_agent_m0_write),                                       //   input,     width = 1,                         .write
		.uav_waitrequest        (mem0_s1_agent_m0_waitrequest),                                 //  output,     width = 1,                         .waitrequest
		.uav_readdatavalid      (mem0_s1_agent_m0_readdatavalid),                               //  output,     width = 1,                         .readdatavalid
		.uav_byteenable         (mem0_s1_agent_m0_byteenable),                                  //   input,   width = 128,                         .byteenable
		.uav_readdata           (mem0_s1_agent_m0_readdata),                                    //  output,  width = 1024,                         .readdata
		.uav_writedata          (mem0_s1_agent_m0_writedata),                                   //   input,  width = 1024,                         .writedata
		.uav_lock               (mem0_s1_agent_m0_lock),                                        //   input,     width = 1,                         .lock
		.uav_debugaccess        (mem0_s1_agent_m0_debugaccess),                                 //   input,     width = 1,                         .debugaccess
		.av_address             (MEM0_s1_address),                                              //  output,     width = 8,      avalon_anti_slave_0.address
		.av_write               (MEM0_s1_write),                                                //  output,     width = 1,                         .write
		.av_readdata            (MEM0_s1_readdata),                                             //   input,  width = 1024,                         .readdata
		.av_writedata           (MEM0_s1_writedata),                                            //  output,  width = 1024,                         .writedata
		.av_byteenable          (MEM0_s1_byteenable),                                           //  output,   width = 128,                         .byteenable
		.av_chipselect          (MEM0_s1_chipselect),                                           //  output,     width = 1,                         .chipselect
		.av_clken               (MEM0_s1_clken),                                                //  output,     width = 1,                         .clken
		.av_read                (),                                                             // (terminated),                                         
		.av_begintransfer       (),                                                             // (terminated),                                         
		.av_beginbursttransfer  (),                                                             // (terminated),                                         
		.av_burstcount          (),                                                             // (terminated),                                         
		.av_readdatavalid       (1'b0),                                                         // (terminated),                                         
		.av_waitrequest         (1'b0),                                                         // (terminated),                                         
		.av_writebyteenable     (),                                                             // (terminated),                                         
		.av_lock                (),                                                             // (terminated),                                         
		.uav_clken              (1'b0),                                                         // (terminated),                                         
		.av_debugaccess         (),                                                             // (terminated),                                         
		.av_outputenable        (),                                                             // (terminated),                                         
		.uav_response           (),                                                             // (terminated),                                         
		.av_response            (2'b00),                                                        // (terminated),                                         
		.uav_writeresponsevalid (),                                                             // (terminated),                                         
		.av_writeresponsevalid  (1'b0)                                                          // (terminated),                                         
	);

	pcie_ed_altera_merlin_master_agent_191_mpbm6tq #(
		.PKT_WUNIQUE               (1266),
		.PKT_DOMAIN_H              (1265),
		.PKT_DOMAIN_L              (1264),
		.PKT_SNOOP_H               (1263),
		.PKT_SNOOP_L               (1260),
		.PKT_BARRIER_H             (1259),
		.PKT_BARRIER_L             (1258),
		.PKT_ORI_BURST_SIZE_H      (1257),
		.PKT_ORI_BURST_SIZE_L      (1255),
		.PKT_RESPONSE_STATUS_H     (1254),
		.PKT_RESPONSE_STATUS_L     (1253),
		.PKT_QOS_H                 (1242),
		.PKT_QOS_L                 (1242),
		.PKT_DATA_SIDEBAND_H       (1240),
		.PKT_DATA_SIDEBAND_L       (1240),
		.PKT_ADDR_SIDEBAND_H       (1239),
		.PKT_ADDR_SIDEBAND_L       (1239),
		.PKT_BURST_TYPE_H          (1238),
		.PKT_BURST_TYPE_L          (1237),
		.PKT_CACHE_H               (1252),
		.PKT_CACHE_L               (1249),
		.PKT_THREAD_ID_H           (1245),
		.PKT_THREAD_ID_L           (1245),
		.PKT_BURST_SIZE_H          (1236),
		.PKT_BURST_SIZE_L          (1234),
		.PKT_TRANS_EXCLUSIVE       (1221),
		.PKT_TRANS_LOCK            (1220),
		.PKT_BEGIN_BURST           (1241),
		.PKT_PROTECTION_H          (1248),
		.PKT_PROTECTION_L          (1246),
		.PKT_BURSTWRAP_H           (1233),
		.PKT_BURSTWRAP_L           (1233),
		.PKT_BYTE_CNT_H            (1232),
		.PKT_BYTE_CNT_L            (1222),
		.PKT_ADDR_H                (1215),
		.PKT_ADDR_L                (1152),
		.PKT_TRANS_COMPRESSED_READ (1216),
		.PKT_TRANS_POSTED          (1217),
		.PKT_TRANS_WRITE           (1218),
		.PKT_TRANS_READ            (1219),
		.PKT_DATA_H                (1023),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (1151),
		.PKT_BYTEEN_L              (1024),
		.PKT_SRC_ID_H              (1243),
		.PKT_SRC_ID_L              (1243),
		.PKT_DEST_ID_H             (1244),
		.PKT_DEST_ID_L             (1244),
		.ST_DATA_W                 (1267),
		.ST_CHANNEL_W              (1),
		.AV_BURSTCOUNT_W           (11),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (1),
		.USE_WRITERESPONSE         (0),
		.DOMAIN_VALUE              (3),
		.BARRIER_VALUE             (0),
		.SNOOP_VALUE               (0),
		.WUNIQUE_VALUE             (0),
		.SYNC_RESET                (1)
	) pio0_pio_master_agent (
		.clk                   (pio0_pio_master_clk_clk),                                            //   input,     width = 1,       clk.clk
		.reset                 (pio0_pio_master_translator_reset_reset_bridge_in_reset_reset),       //   input,     width = 1, clk_reset.reset
		.av_address            (pio0_pio_master_translator_avalon_universal_master_0_address),       //   input,    width = 64,        av.address
		.av_write              (pio0_pio_master_translator_avalon_universal_master_0_write),         //   input,     width = 1,          .write
		.av_read               (pio0_pio_master_translator_avalon_universal_master_0_read),          //   input,     width = 1,          .read
		.av_writedata          (pio0_pio_master_translator_avalon_universal_master_0_writedata),     //   input,  width = 1024,          .writedata
		.av_readdata           (pio0_pio_master_translator_avalon_universal_master_0_readdata),      //  output,  width = 1024,          .readdata
		.av_waitrequest        (pio0_pio_master_translator_avalon_universal_master_0_waitrequest),   //  output,     width = 1,          .waitrequest
		.av_readdatavalid      (pio0_pio_master_translator_avalon_universal_master_0_readdatavalid), //  output,     width = 1,          .readdatavalid
		.av_byteenable         (pio0_pio_master_translator_avalon_universal_master_0_byteenable),    //   input,   width = 128,          .byteenable
		.av_burstcount         (pio0_pio_master_translator_avalon_universal_master_0_burstcount),    //   input,    width = 11,          .burstcount
		.av_debugaccess        (pio0_pio_master_translator_avalon_universal_master_0_debugaccess),   //   input,     width = 1,          .debugaccess
		.av_lock               (pio0_pio_master_translator_avalon_universal_master_0_lock),          //   input,     width = 1,          .lock
		.av_response           (pio0_pio_master_translator_avalon_universal_master_0_response),      //  output,     width = 2,          .response
		.cp_valid              (pio0_pio_master_agent_cp_valid),                                     //  output,     width = 1,        cp.valid
		.cp_data               (pio0_pio_master_agent_cp_data),                                      //  output,  width = 1267,          .data
		.cp_startofpacket      (pio0_pio_master_agent_cp_startofpacket),                             //  output,     width = 1,          .startofpacket
		.cp_endofpacket        (pio0_pio_master_agent_cp_endofpacket),                               //  output,     width = 1,          .endofpacket
		.cp_ready              (pio0_pio_master_agent_cp_ready),                                     //   input,     width = 1,          .ready
		.rp_valid              (rsp_mux_src_valid),                                                  //   input,     width = 1,        rp.valid
		.rp_data               (rsp_mux_src_data),                                                   //   input,  width = 1267,          .data
		.rp_channel            (rsp_mux_src_channel),                                                //   input,     width = 1,          .channel
		.rp_startofpacket      (rsp_mux_src_startofpacket),                                          //   input,     width = 1,          .startofpacket
		.rp_endofpacket        (rsp_mux_src_endofpacket),                                            //   input,     width = 1,          .endofpacket
		.rp_ready              (rsp_mux_src_ready),                                                  //  output,     width = 1,          .ready
		.av_writeresponsevalid ()                                                                    // (terminated),                          
	);

	pcie_ed_altera_merlin_slave_agent_191_ncfkfri #(
		.PKT_ORI_BURST_SIZE_H      (1257),
		.PKT_ORI_BURST_SIZE_L      (1255),
		.PKT_RESPONSE_STATUS_H     (1254),
		.PKT_RESPONSE_STATUS_L     (1253),
		.PKT_BURST_SIZE_H          (1236),
		.PKT_BURST_SIZE_L          (1234),
		.PKT_TRANS_LOCK            (1220),
		.PKT_BEGIN_BURST           (1241),
		.PKT_PROTECTION_H          (1248),
		.PKT_PROTECTION_L          (1246),
		.PKT_BURSTWRAP_H           (1233),
		.PKT_BURSTWRAP_L           (1233),
		.PKT_BYTE_CNT_H            (1232),
		.PKT_BYTE_CNT_L            (1222),
		.PKT_ADDR_H                (1215),
		.PKT_ADDR_L                (1152),
		.PKT_TRANS_COMPRESSED_READ (1216),
		.PKT_TRANS_POSTED          (1217),
		.PKT_TRANS_WRITE           (1218),
		.PKT_TRANS_READ            (1219),
		.PKT_DATA_H                (1023),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (1151),
		.PKT_BYTEEN_L              (1024),
		.PKT_SRC_ID_H              (1243),
		.PKT_SRC_ID_L              (1243),
		.PKT_DEST_ID_H             (1244),
		.PKT_DEST_ID_L             (1244),
		.PKT_SYMBOL_W              (8),
		.ST_CHANNEL_W              (1),
		.ST_DATA_W                 (1267),
		.AVS_BURSTCOUNT_W          (8),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0),
		.ECC_ENABLE                (0),
		.SYNC_RESET                (1)
	) mem0_s1_agent (
		.clk                     (pio0_pio_master_clk_clk),                                      //   input,     width = 1,             clk.clk
		.reset                   (pio0_pio_master_translator_reset_reset_bridge_in_reset_reset), //   input,     width = 1,       clk_reset.reset
		.m0_address              (mem0_s1_agent_m0_address),                                     //  output,    width = 64,              m0.address
		.m0_burstcount           (mem0_s1_agent_m0_burstcount),                                  //  output,     width = 8,                .burstcount
		.m0_byteenable           (mem0_s1_agent_m0_byteenable),                                  //  output,   width = 128,                .byteenable
		.m0_debugaccess          (mem0_s1_agent_m0_debugaccess),                                 //  output,     width = 1,                .debugaccess
		.m0_lock                 (mem0_s1_agent_m0_lock),                                        //  output,     width = 1,                .lock
		.m0_readdata             (mem0_s1_agent_m0_readdata),                                    //   input,  width = 1024,                .readdata
		.m0_readdatavalid        (mem0_s1_agent_m0_readdatavalid),                               //   input,     width = 1,                .readdatavalid
		.m0_read                 (mem0_s1_agent_m0_read),                                        //  output,     width = 1,                .read
		.m0_waitrequest          (mem0_s1_agent_m0_waitrequest),                                 //   input,     width = 1,                .waitrequest
		.m0_writedata            (mem0_s1_agent_m0_writedata),                                   //  output,  width = 1024,                .writedata
		.m0_write                (mem0_s1_agent_m0_write),                                       //  output,     width = 1,                .write
		.rp_endofpacket          (mem0_s1_agent_rp_endofpacket),                                 //  output,     width = 1,              rp.endofpacket
		.rp_ready                (mem0_s1_agent_rp_ready),                                       //   input,     width = 1,                .ready
		.rp_valid                (mem0_s1_agent_rp_valid),                                       //  output,     width = 1,                .valid
		.rp_data                 (mem0_s1_agent_rp_data),                                        //  output,  width = 1267,                .data
		.rp_startofpacket        (mem0_s1_agent_rp_startofpacket),                               //  output,     width = 1,                .startofpacket
		.cp_ready                (mem0_s1_burst_adapter_source0_ready),                          //  output,     width = 1,              cp.ready
		.cp_valid                (mem0_s1_burst_adapter_source0_valid),                          //   input,     width = 1,                .valid
		.cp_data                 (mem0_s1_burst_adapter_source0_data),                           //   input,  width = 1267,                .data
		.cp_startofpacket        (mem0_s1_burst_adapter_source0_startofpacket),                  //   input,     width = 1,                .startofpacket
		.cp_endofpacket          (mem0_s1_burst_adapter_source0_endofpacket),                    //   input,     width = 1,                .endofpacket
		.cp_channel              (mem0_s1_burst_adapter_source0_channel),                        //   input,     width = 1,                .channel
		.rf_sink_ready           (mem0_s1_agent_rsp_fifo_out_ready),                             //  output,     width = 1,         rf_sink.ready
		.rf_sink_valid           (mem0_s1_agent_rsp_fifo_out_valid),                             //   input,     width = 1,                .valid
		.rf_sink_startofpacket   (mem0_s1_agent_rsp_fifo_out_startofpacket),                     //   input,     width = 1,                .startofpacket
		.rf_sink_endofpacket     (mem0_s1_agent_rsp_fifo_out_endofpacket),                       //   input,     width = 1,                .endofpacket
		.rf_sink_data            (mem0_s1_agent_rsp_fifo_out_data),                              //   input,  width = 1268,                .data
		.rf_source_ready         (mem0_s1_agent_rf_source_ready),                                //   input,     width = 1,       rf_source.ready
		.rf_source_valid         (mem0_s1_agent_rf_source_valid),                                //  output,     width = 1,                .valid
		.rf_source_startofpacket (mem0_s1_agent_rf_source_startofpacket),                        //  output,     width = 1,                .startofpacket
		.rf_source_endofpacket   (mem0_s1_agent_rf_source_endofpacket),                          //  output,     width = 1,                .endofpacket
		.rf_source_data          (mem0_s1_agent_rf_source_data),                                 //  output,  width = 1268,                .data
		.rdata_fifo_sink_ready   (mem0_s1_agent_rdata_fifo_src_ready),                           //  output,     width = 1, rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (mem0_s1_agent_rdata_fifo_src_valid),                           //   input,     width = 1,                .valid
		.rdata_fifo_sink_data    (mem0_s1_agent_rdata_fifo_src_data),                            //   input,  width = 1026,                .data
		.rdata_fifo_src_ready    (mem0_s1_agent_rdata_fifo_src_ready),                           //   input,     width = 1,  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (mem0_s1_agent_rdata_fifo_src_valid),                           //  output,     width = 1,                .valid
		.rdata_fifo_src_data     (mem0_s1_agent_rdata_fifo_src_data),                            //  output,  width = 1026,                .data
		.m0_response             (2'b00),                                                        // (terminated),                                
		.m0_writeresponsevalid   (1'b0),                                                         // (terminated),                                
		.rdata_fifo_sink_error   (1'b0)                                                          // (terminated),                                
	);

	pcie_ed_altera_avalon_sc_fifo_1931_vhmcgqy #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (1268),
		.FIFO_DEPTH          (3),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0),
		.EMPTY_WIDTH         (1),
		.SYNC_RESET          (1)
	) mem0_s1_agent_rsp_fifo (
		.clk               (pio0_pio_master_clk_clk),                  //   input,     width = 1,       clk.clk
		.reset             (MEM0_reset1_reset_bridge_in_reset_reset),  //   input,     width = 1, clk_reset.reset
		.in_data           (mem0_s1_agent_rf_source_data),             //   input,  width = 1268,        in.data
		.in_valid          (mem0_s1_agent_rf_source_valid),            //   input,     width = 1,          .valid
		.in_ready          (mem0_s1_agent_rf_source_ready),            //  output,     width = 1,          .ready
		.in_startofpacket  (mem0_s1_agent_rf_source_startofpacket),    //   input,     width = 1,          .startofpacket
		.in_endofpacket    (mem0_s1_agent_rf_source_endofpacket),      //   input,     width = 1,          .endofpacket
		.out_data          (mem0_s1_agent_rsp_fifo_out_data),          //  output,  width = 1268,       out.data
		.out_valid         (mem0_s1_agent_rsp_fifo_out_valid),         //  output,     width = 1,          .valid
		.out_ready         (mem0_s1_agent_rsp_fifo_out_ready),         //   input,     width = 1,          .ready
		.out_startofpacket (mem0_s1_agent_rsp_fifo_out_startofpacket), //  output,     width = 1,          .startofpacket
		.out_endofpacket   (mem0_s1_agent_rsp_fifo_out_endofpacket),   //  output,     width = 1,          .endofpacket
		.csr_address       (2'b00),                                    // (terminated),                          
		.csr_read          (1'b0),                                     // (terminated),                          
		.csr_write         (1'b0),                                     // (terminated),                          
		.csr_readdata      (),                                         // (terminated),                          
		.csr_writedata     (32'b00000000000000000000000000000000),     // (terminated),                          
		.almost_full_data  (),                                         // (terminated),                          
		.almost_empty_data (),                                         // (terminated),                          
		.in_empty          (1'b0),                                     // (terminated),                          
		.out_empty         (),                                         // (terminated),                          
		.in_error          (1'b0),                                     // (terminated),                          
		.out_error         (),                                         // (terminated),                          
		.in_channel        (1'b0),                                     // (terminated),                          
		.out_channel       ()                                          // (terminated),                          
	);

	pcie_ed_altera_merlin_router_1921_6kkcoeq router (
		.sink_ready         (pio0_pio_master_agent_cp_ready),                               //  output,     width = 1,      sink.ready
		.sink_valid         (pio0_pio_master_agent_cp_valid),                               //   input,     width = 1,          .valid
		.sink_data          (pio0_pio_master_agent_cp_data),                                //   input,  width = 1267,          .data
		.sink_startofpacket (pio0_pio_master_agent_cp_startofpacket),                       //   input,     width = 1,          .startofpacket
		.sink_endofpacket   (pio0_pio_master_agent_cp_endofpacket),                         //   input,     width = 1,          .endofpacket
		.clk                (pio0_pio_master_clk_clk),                                      //   input,     width = 1,       clk.clk
		.reset              (pio0_pio_master_translator_reset_reset_bridge_in_reset_reset), //   input,     width = 1, clk_reset.reset
		.src_ready          (router_src_ready),                                             //   input,     width = 1,       src.ready
		.src_valid          (router_src_valid),                                             //  output,     width = 1,          .valid
		.src_data           (router_src_data),                                              //  output,  width = 1267,          .data
		.src_channel        (router_src_channel),                                           //  output,     width = 1,          .channel
		.src_startofpacket  (router_src_startofpacket),                                     //  output,     width = 1,          .startofpacket
		.src_endofpacket    (router_src_endofpacket)                                        //  output,     width = 1,          .endofpacket
	);

	pcie_ed_altera_merlin_router_1921_sv2vwxi router_001 (
		.sink_ready         (mem0_s1_agent_rp_ready),                                       //  output,     width = 1,      sink.ready
		.sink_valid         (mem0_s1_agent_rp_valid),                                       //   input,     width = 1,          .valid
		.sink_data          (mem0_s1_agent_rp_data),                                        //   input,  width = 1267,          .data
		.sink_startofpacket (mem0_s1_agent_rp_startofpacket),                               //   input,     width = 1,          .startofpacket
		.sink_endofpacket   (mem0_s1_agent_rp_endofpacket),                                 //   input,     width = 1,          .endofpacket
		.clk                (pio0_pio_master_clk_clk),                                      //   input,     width = 1,       clk.clk
		.reset              (pio0_pio_master_translator_reset_reset_bridge_in_reset_reset), //   input,     width = 1, clk_reset.reset
		.src_ready          (router_001_src_ready),                                         //   input,     width = 1,       src.ready
		.src_valid          (router_001_src_valid),                                         //  output,     width = 1,          .valid
		.src_data           (router_001_src_data),                                          //  output,  width = 1267,          .data
		.src_channel        (router_001_src_channel),                                       //  output,     width = 1,          .channel
		.src_startofpacket  (router_001_src_startofpacket),                                 //  output,     width = 1,          .startofpacket
		.src_endofpacket    (router_001_src_endofpacket)                                    //  output,     width = 1,          .endofpacket
	);

	pcie_ed_altera_merlin_burst_adapter_1922_tsepz7q #(
		.PKT_ADDR_H                (1215),
		.PKT_ADDR_L                (1152),
		.PKT_BEGIN_BURST           (1241),
		.PKT_BYTE_CNT_H            (1232),
		.PKT_BYTE_CNT_L            (1222),
		.PKT_BYTEEN_H              (1151),
		.PKT_BYTEEN_L              (1024),
		.PKT_BURST_SIZE_H          (1236),
		.PKT_BURST_SIZE_L          (1234),
		.PKT_BURST_TYPE_H          (1238),
		.PKT_BURST_TYPE_L          (1237),
		.PKT_BURSTWRAP_H           (1233),
		.PKT_BURSTWRAP_L           (1233),
		.PKT_TRANS_COMPRESSED_READ (1216),
		.PKT_TRANS_WRITE           (1218),
		.PKT_TRANS_READ            (1219),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (1267),
		.ST_CHANNEL_W              (1),
		.OUT_BYTE_CNT_H            (1229),
		.OUT_BURSTWRAP_H           (1233),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.INCOMPLETE_WRAP_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (1),
		.BURSTWRAP_CONST_VALUE     (1),
		.ADAPTER_VERSION           ("13.1"),
		.SYNC_RESET                (1)
	) mem0_s1_burst_adapter (
		.clk                   (pio0_pio_master_clk_clk),                                      //   input,     width = 1,       cr0.clk
		.reset                 (pio0_pio_master_translator_reset_reset_bridge_in_reset_reset), //   input,     width = 1, cr0_reset.reset
		.sink0_valid           (cmd_mux_src_valid),                                            //   input,     width = 1,     sink0.valid
		.sink0_data            (cmd_mux_src_data),                                             //   input,  width = 1267,          .data
		.sink0_channel         (cmd_mux_src_channel),                                          //   input,     width = 1,          .channel
		.sink0_startofpacket   (cmd_mux_src_startofpacket),                                    //   input,     width = 1,          .startofpacket
		.sink0_endofpacket     (cmd_mux_src_endofpacket),                                      //   input,     width = 1,          .endofpacket
		.sink0_ready           (cmd_mux_src_ready),                                            //  output,     width = 1,          .ready
		.source0_valid         (mem0_s1_burst_adapter_source0_valid),                          //  output,     width = 1,   source0.valid
		.source0_data          (mem0_s1_burst_adapter_source0_data),                           //  output,  width = 1267,          .data
		.source0_channel       (mem0_s1_burst_adapter_source0_channel),                        //  output,     width = 1,          .channel
		.source0_startofpacket (mem0_s1_burst_adapter_source0_startofpacket),                  //  output,     width = 1,          .startofpacket
		.source0_endofpacket   (mem0_s1_burst_adapter_source0_endofpacket),                    //  output,     width = 1,          .endofpacket
		.source0_ready         (mem0_s1_burst_adapter_source0_ready)                           //   input,     width = 1,          .ready
	);

	pcie_ed_altera_merlin_demultiplexer_1921_s5kn7vi cmd_demux (
		.clk                (pio0_pio_master_clk_clk),                                      //   input,     width = 1,       clk.clk
		.reset              (pio0_pio_master_translator_reset_reset_bridge_in_reset_reset), //   input,     width = 1, clk_reset.reset
		.sink_ready         (router_src_ready),                                             //  output,     width = 1,      sink.ready
		.sink_channel       (router_src_channel),                                           //   input,     width = 1,          .channel
		.sink_data          (router_src_data),                                              //   input,  width = 1267,          .data
		.sink_startofpacket (router_src_startofpacket),                                     //   input,     width = 1,          .startofpacket
		.sink_endofpacket   (router_src_endofpacket),                                       //   input,     width = 1,          .endofpacket
		.sink_valid         (router_src_valid),                                             //   input,     width = 1,          .valid
		.src0_ready         (cmd_demux_src0_ready),                                         //   input,     width = 1,      src0.ready
		.src0_valid         (cmd_demux_src0_valid),                                         //  output,     width = 1,          .valid
		.src0_data          (cmd_demux_src0_data),                                          //  output,  width = 1267,          .data
		.src0_channel       (cmd_demux_src0_channel),                                       //  output,     width = 1,          .channel
		.src0_startofpacket (cmd_demux_src0_startofpacket),                                 //  output,     width = 1,          .startofpacket
		.src0_endofpacket   (cmd_demux_src0_endofpacket)                                    //  output,     width = 1,          .endofpacket
	);

	pcie_ed_altera_merlin_multiplexer_1921_zxmqgaq cmd_mux (
		.clk                 (pio0_pio_master_clk_clk),                                      //   input,     width = 1,       clk.clk
		.reset               (pio0_pio_master_translator_reset_reset_bridge_in_reset_reset), //   input,     width = 1, clk_reset.reset
		.src_ready           (cmd_mux_src_ready),                                            //   input,     width = 1,       src.ready
		.src_valid           (cmd_mux_src_valid),                                            //  output,     width = 1,          .valid
		.src_data            (cmd_mux_src_data),                                             //  output,  width = 1267,          .data
		.src_channel         (cmd_mux_src_channel),                                          //  output,     width = 1,          .channel
		.src_startofpacket   (cmd_mux_src_startofpacket),                                    //  output,     width = 1,          .startofpacket
		.src_endofpacket     (cmd_mux_src_endofpacket),                                      //  output,     width = 1,          .endofpacket
		.sink0_ready         (cmd_demux_src0_ready),                                         //  output,     width = 1,     sink0.ready
		.sink0_valid         (cmd_demux_src0_valid),                                         //   input,     width = 1,          .valid
		.sink0_channel       (cmd_demux_src0_channel),                                       //   input,     width = 1,          .channel
		.sink0_data          (cmd_demux_src0_data),                                          //   input,  width = 1267,          .data
		.sink0_startofpacket (cmd_demux_src0_startofpacket),                                 //   input,     width = 1,          .startofpacket
		.sink0_endofpacket   (cmd_demux_src0_endofpacket)                                    //   input,     width = 1,          .endofpacket
	);

	pcie_ed_altera_merlin_demultiplexer_1921_s5kn7vi rsp_demux (
		.clk                (pio0_pio_master_clk_clk),                                      //   input,     width = 1,       clk.clk
		.reset              (pio0_pio_master_translator_reset_reset_bridge_in_reset_reset), //   input,     width = 1, clk_reset.reset
		.sink_ready         (router_001_src_ready),                                         //  output,     width = 1,      sink.ready
		.sink_channel       (router_001_src_channel),                                       //   input,     width = 1,          .channel
		.sink_data          (router_001_src_data),                                          //   input,  width = 1267,          .data
		.sink_startofpacket (router_001_src_startofpacket),                                 //   input,     width = 1,          .startofpacket
		.sink_endofpacket   (router_001_src_endofpacket),                                   //   input,     width = 1,          .endofpacket
		.sink_valid         (router_001_src_valid),                                         //   input,     width = 1,          .valid
		.src0_ready         (rsp_demux_src0_ready),                                         //   input,     width = 1,      src0.ready
		.src0_valid         (rsp_demux_src0_valid),                                         //  output,     width = 1,          .valid
		.src0_data          (rsp_demux_src0_data),                                          //  output,  width = 1267,          .data
		.src0_channel       (rsp_demux_src0_channel),                                       //  output,     width = 1,          .channel
		.src0_startofpacket (rsp_demux_src0_startofpacket),                                 //  output,     width = 1,          .startofpacket
		.src0_endofpacket   (rsp_demux_src0_endofpacket)                                    //  output,     width = 1,          .endofpacket
	);

	pcie_ed_altera_merlin_multiplexer_1921_5zcdh2i rsp_mux (
		.clk                 (pio0_pio_master_clk_clk),                                      //   input,     width = 1,       clk.clk
		.reset               (pio0_pio_master_translator_reset_reset_bridge_in_reset_reset), //   input,     width = 1, clk_reset.reset
		.src_ready           (rsp_mux_src_ready),                                            //   input,     width = 1,       src.ready
		.src_valid           (rsp_mux_src_valid),                                            //  output,     width = 1,          .valid
		.src_data            (rsp_mux_src_data),                                             //  output,  width = 1267,          .data
		.src_channel         (rsp_mux_src_channel),                                          //  output,     width = 1,          .channel
		.src_startofpacket   (rsp_mux_src_startofpacket),                                    //  output,     width = 1,          .startofpacket
		.src_endofpacket     (rsp_mux_src_endofpacket),                                      //  output,     width = 1,          .endofpacket
		.sink0_ready         (rsp_demux_src0_ready),                                         //  output,     width = 1,     sink0.ready
		.sink0_valid         (rsp_demux_src0_valid),                                         //   input,     width = 1,          .valid
		.sink0_channel       (rsp_demux_src0_channel),                                       //   input,     width = 1,          .channel
		.sink0_data          (rsp_demux_src0_data),                                          //   input,  width = 1267,          .data
		.sink0_startofpacket (rsp_demux_src0_startofpacket),                                 //   input,     width = 1,          .startofpacket
		.sink0_endofpacket   (rsp_demux_src0_endofpacket)                                    //   input,     width = 1,          .endofpacket
	);

endmodule
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "EtAh8aN7m2BPKOTfO5tEAbNSD19BnNEklF4xQRY7YZ2oRe/8wDIRx8XCKuwkXQtjYcM5gRXSD6c+oGX77mfnvlAGw9KTmnXPBu3GU7e3qFjUTrXWlEAN76gMqJTePk91Iv2qtpAKuY2LJHLiowUVDoSuAt1Csh1O2u7qDzQRIaeVL/AJWYDMfWERE2K26wZcHHB8eTbMnhSND4m01aQODfKXixyUFYBUVJCy/gZrUwDQOCgsvIWE/ANcrGEWYMvIzvknETHHBWq7hvzRDCTNQp32gjZBXno1lGnDCN9nhYslMrOhArI8PPAgnnT3gDwF0Kc6Ef2kybQo7er/WTqXu0imPKaM5V5eGwkLxZlEAlTUKTBb4lV3MK7fLUvRplvQHXx9VlEtifqdLc6rPX5czWFPomkKm1K+w0jx8/msm9sX8LEEt+2get+E0Z91Vj6Ltj7Gc+FCqKufoYvp6mLFdkDBOfizPwrJ9Z1PPd5AetIWoxKltH6vnAKlCndphzV9wLTpdimgIJnO07ljzzawk9uoiGRWX5uYqNZgX+92d2nfsawrGO0BQaj5K/2za6KYFHKwNDYbyuv4K1FyJO2t9eTNEqt1VN51uf2tTqzTm6HjoaIq/6DYepMghg35wfuI4Li2fgoxB6dlov4U1F4OgyxrjJ6jxhgah4iPR6GCnOqgGJ4e9ZLlrbfLG1rFRro/O6uvuzTOl9uSpuMRoV04J7pGq6ALlwUVXXjpkOTV5LVBHjoGGE2y7QhKkLS2ziDk5fZHMk6M4cuhK1lOa2fL6wAxU3J4lO7QBNxa40qljvbMlYkwv32UHWLV+xjgJfiR8jmKXpDLwADkAS4EoTYmFbjVQHuseb8/8ZEGnGFDluS7z7Wg3MR/LndSC1VUlZUM1Kj8adFzOZ7rswL/I9wBcWJQxh+gaQAvfGzq/FePg48fhhvGEO8YYHV/2jNDQaeZgqIuwvKtMvR9+tI7bnQaZjUKaYfTeUljNMp4l3HEZ6Sqadjk5Hpk+c/YsvysDd2Z"
`endif